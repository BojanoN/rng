/* Verilog model created from schematic x.sch -- Jan 21, 2016 23:35 */

module x;



OB I1 ();

endmodule // x
